module left_shift_32 (res, data, select);
input[31:0] data;
input[4:0] select;
output[31:0] res;
wire[31:0] W1, W2, W3, W4;  //intermediate carries
// mux_2_1_helper(result, d, s)

//LEVEL 1 SHIFT
mux_2_1_helper mux0(W1[0], 1'b0 , data[0], select[0]);
mux_2_1_helper mux1(W1[1], data[0] , data[1], select[0]);
mux_2_1_helper mux2(W1[2], data[1] , data[2], select[0]);
mux_2_1_helper mux3(W1[3], data[2] , data[3], select[0]);
mux_2_1_helper mux4(W1[4], data[3] , data[4], select[0]);
mux_2_1_helper mux5(W1[5], data[4] , data[5], select[0]);
mux_2_1_helper mux6(W1[6], data[5] , data[6], select[0]);
mux_2_1_helper mux7(W1[7], data[6] , data[7], select[0]);
mux_2_1_helper mux8(W1[8], data[7] , data[8], select[0]);
mux_2_1_helper mux9(W1[9], data[8] , data[9], select[0]);
mux_2_1_helper mux10(W1[10], data[9] , data[10], select[0]);
mux_2_1_helper mux11(W1[11], data[10] , data[11], select[0]);
mux_2_1_helper mux12(W1[12], data[11] , data[12], select[0]);
mux_2_1_helper mux13(W1[13], data[12] , data[13], select[0]);
mux_2_1_helper mux14(W1[14], data[13] , data[14], select[0]);
mux_2_1_helper mux15(W1[15], data[14] , data[15], select[0]);
mux_2_1_helper mux16(W1[16], data[15] , data[16], select[0]);
mux_2_1_helper mux17(W1[17], data[16] , data[17], select[0]);
mux_2_1_helper mux18(W1[18], data[17] , data[18], select[0]);
mux_2_1_helper mux19(W1[19], data[18] , data[19], select[0]);
mux_2_1_helper mux20(W1[20], data[19] , data[20], select[0]);
mux_2_1_helper mux21(W1[21], data[20] , data[21], select[0]);
mux_2_1_helper mux22(W1[22], data[21] , data[22], select[0]);
mux_2_1_helper mux23(W1[23], data[22] , data[23], select[0]);
mux_2_1_helper mux24(W1[24], data[23] , data[24], select[0]);
mux_2_1_helper mux25(W1[25], data[24] , data[25], select[0]);
mux_2_1_helper mux26(W1[26], data[25] , data[26], select[0]);
mux_2_1_helper mux27(W1[27], data[26] , data[27], select[0]);
mux_2_1_helper mux28(W1[28], data[27] , data[28], select[0]);
mux_2_1_helper mux29(W1[29], data[28] , data[29], select[0]);
mux_2_1_helper mux30(W1[30], data[29] , data[30], select[0]);
mux_2_1_helper mux31(W1[31], data[30] , data[31], select[0]);

//LEVEL 2 SHIFT
mux_2_1_helper mux33(W2[0], 1'b0 , W1[0], select[1]);
mux_2_1_helper mux34(W2[1], 1'b0 , W1[1], select[1]);
mux_2_1_helper mux35(W2[2], W1[0] , W1[2], select[1]);
mux_2_1_helper mux36(W2[3], W1[1] , W1[3], select[1]);
mux_2_1_helper mux37(W2[4], W1[2] , W1[4], select[1]);
mux_2_1_helper mux38(W2[5], W1[3] , W1[5], select[1]);
mux_2_1_helper mux39(W2[6], W1[4] , W1[6], select[1]);
mux_2_1_helper mux40(W2[7], W1[5] , W1[7], select[1]);
mux_2_1_helper mux41(W2[8], W1[6] , W1[8], select[1]);
mux_2_1_helper mux42(W2[9], W1[7] , W1[9], select[1]);
mux_2_1_helper mux43(W2[10], W1[8] , W1[10], select[1]);
mux_2_1_helper mux44(W2[11], W1[9] , W1[11], select[1]);
mux_2_1_helper mux45(W2[12], W1[10] , W1[12], select[1]);
mux_2_1_helper mux46(W2[13], W1[11] , W1[13], select[1]);
mux_2_1_helper mux47(W2[14], W1[12] , W1[14], select[1]);
mux_2_1_helper mux48(W2[15], W1[13] , W1[15], select[1]);
mux_2_1_helper mux49(W2[16], W1[14] , W1[16], select[1]);
mux_2_1_helper mux50(W2[17], W1[15] , W1[17], select[1]);
mux_2_1_helper mux51(W2[18], W1[16] , W1[18], select[1]);
mux_2_1_helper mux52(W2[19], W1[17] , W1[19], select[1]);
mux_2_1_helper mux53(W2[20], W1[18] , W1[20], select[1]);
mux_2_1_helper mux54(W2[21], W1[19] , W1[21], select[1]);
mux_2_1_helper mux55(W2[22], W1[20] , W1[22], select[1]);
mux_2_1_helper mux56(W2[23], W1[21] , W1[23], select[1]);
mux_2_1_helper mux57(W2[24], W1[22] , W1[24], select[1]);
mux_2_1_helper mux58(W2[25], W1[23] , W1[25], select[1]);
mux_2_1_helper mux59(W2[26], W1[24] , W1[26], select[1]);
mux_2_1_helper mux60(W2[27], W1[25] , W1[27], select[1]);
mux_2_1_helper mux61(W2[28], W1[26] , W1[28], select[1]);
mux_2_1_helper mux62(W2[29], W1[27] , W1[29], select[1]);
mux_2_1_helper mux63(W2[30], W1[28] , W1[30], select[1]);
mux_2_1_helper mux64(W2[31], W1[29] , W1[31], select[1]);

//LEVEL 3 SHIFT
mux_2_1_helper mux65(W3[0], 1'b0 , W2[0], select[2]);
mux_2_1_helper mux66(W3[1], 1'b0 , W2[1], select[2]);
mux_2_1_helper mux67(W3[2], 1'b0 , W2[2], select[2]);
mux_2_1_helper mux68(W3[3], 1'b0 , W2[3], select[2]);
mux_2_1_helper mux69(W3[4], W2[0] , W2[4], select[2]);
mux_2_1_helper mux70(W3[5], W2[1] , W2[5], select[2]);
mux_2_1_helper mux71(W3[6], W2[2] , W2[6], select[2]);
mux_2_1_helper mux72(W3[7], W2[3] , W2[7], select[2]);
mux_2_1_helper mux73(W3[8], W2[4] , W2[8], select[2]);
mux_2_1_helper mux74(W3[9], W2[5] , W2[9], select[2]);
mux_2_1_helper mux75(W3[10], W2[6] , W2[10], select[2]);
mux_2_1_helper mux76(W3[11], W2[7] , W2[11], select[2]);
mux_2_1_helper mux77(W3[12], W2[8] , W2[12], select[2]);
mux_2_1_helper mux78(W3[13], W2[9] , W2[13], select[2]);
mux_2_1_helper mux79(W3[14], W2[10] , W2[14], select[2]);
mux_2_1_helper mux80(W3[15], W2[11] , W2[15], select[2]);
mux_2_1_helper mux81(W3[16], W2[12] , W2[16], select[2]);
mux_2_1_helper mux82(W3[17], W2[13] , W2[17], select[2]);
mux_2_1_helper mux83(W3[18], W2[14] , W2[18], select[2]);
mux_2_1_helper mux84(W3[19], W2[15] , W2[19], select[2]);
mux_2_1_helper mux85(W3[20], W2[16] , W2[20], select[2]);
mux_2_1_helper mux86(W3[21], W2[17] , W2[21], select[2]);
mux_2_1_helper mux87(W3[22], W2[18] , W2[22], select[2]);
mux_2_1_helper mux88(W3[23], W2[19] , W2[23], select[2]);
mux_2_1_helper mux89(W3[24], W2[20] , W2[24], select[2]);
mux_2_1_helper mux90(W3[25], W2[21] , W2[25], select[2]);
mux_2_1_helper mux91(W3[26], W2[22] , W2[26], select[2]);
mux_2_1_helper mux92(W3[27], W2[23] , W2[27], select[2]);
mux_2_1_helper mux93(W3[28], W2[24] , W2[28], select[2]);
mux_2_1_helper mux94(W3[29], W2[25] , W2[29], select[2]);
mux_2_1_helper mux95(W3[30], W2[26] , W2[30], select[2]);
mux_2_1_helper mux96(W3[31], W2[27] , W2[31], select[2]);

//LEVEL 4 SHIFT
mux_2_1_helper mux97(W4[0], 1'b0 , W3[0], select[3]);
mux_2_1_helper mux98(W4[1], 1'b0 , W3[1], select[3]);
mux_2_1_helper mux99(W4[2], 1'b0 , W3[2], select[3]);
mux_2_1_helper mux100(W4[3], 1'b0 , W3[3], select[3]);
mux_2_1_helper mux101(W4[4], 1'b0 , W3[4], select[3]);
mux_2_1_helper mux102(W4[5], 1'b0 , W3[5], select[3]);
mux_2_1_helper mux103(W4[6], 1'b0 , W3[6], select[3]);
mux_2_1_helper mux104(W4[7], 1'b0 , W3[7], select[3]);
mux_2_1_helper mux105(W4[8], W3[0] , W3[8], select[3]);
mux_2_1_helper mux106(W4[9], W3[1] , W3[9], select[3]);
mux_2_1_helper mux107(W4[10], W3[2] , W3[10], select[3]);
mux_2_1_helper mux108(W4[11], W3[3] , W3[11], select[3]);
mux_2_1_helper mux109(W4[12], W3[4] , W3[12], select[3]);
mux_2_1_helper mux110(W4[13], W3[5] , W3[13], select[3]);
mux_2_1_helper mux111(W4[14], W3[6] , W3[14], select[3]);
mux_2_1_helper mux112(W4[15], W3[7] , W3[15], select[3]);
mux_2_1_helper mux113(W4[16], W3[8] , W3[16], select[3]);
mux_2_1_helper mux114(W4[17], W3[9] , W3[17], select[3]);
mux_2_1_helper mux115(W4[18], W3[10] , W3[18], select[3]);
mux_2_1_helper mux116(W4[19], W3[11] , W3[19], select[3]);
mux_2_1_helper mux117(W4[20], W3[12] , W3[20], select[3]);
mux_2_1_helper mux118(W4[21], W3[13] , W3[21], select[3]);
mux_2_1_helper mux119(W4[22], W3[14] , W3[22], select[3]);
mux_2_1_helper mux120(W4[23], W3[15] , W3[23], select[3]);
mux_2_1_helper mux121(W4[24], W3[16] , W3[24], select[3]);
mux_2_1_helper mux122(W4[25], W3[17] , W3[25], select[3]);
mux_2_1_helper mux123(W4[26], W3[18] , W3[26], select[3]);
mux_2_1_helper mux124(W4[27], W3[19] , W3[27], select[3]);
mux_2_1_helper mux125(W4[28], W3[20] , W3[28], select[3]);
mux_2_1_helper mux126(W4[29], W3[21] , W3[29], select[3]);
mux_2_1_helper mux127(W4[30], W3[22] , W3[30], select[3]);
mux_2_1_helper mux128(W4[31], W3[23] , W3[31], select[3]);

//LEVEL 5 SHIFT
mux_2_1_helper mux129(res[0], 1'b0 , W4[0], select[4]);
mux_2_1_helper mux130(res[1], 1'b0 , W4[1], select[4]);
mux_2_1_helper mux131(res[2], 1'b0 , W4[2], select[4]);
mux_2_1_helper mux132(res[3], 1'b0 , W4[3], select[4]);
mux_2_1_helper mux133(res[4], 1'b0 , W4[4], select[4]);
mux_2_1_helper mux134(res[5], 1'b0 , W4[5], select[4]);
mux_2_1_helper mux135(res[6], 1'b0 , W4[6], select[4]);
mux_2_1_helper mux136(res[7], 1'b0 , W4[7], select[4]);
mux_2_1_helper mux137(res[8], 1'b0 , W4[8], select[4]);
mux_2_1_helper mux138(res[9], 1'b0 , W4[9], select[4]);
mux_2_1_helper mux139(res[10], 1'b0 , W4[10], select[4]);
mux_2_1_helper mux140(res[11], 1'b0 , W4[11], select[4]);
mux_2_1_helper mux141(res[12], 1'b0 , W4[12], select[4]);
mux_2_1_helper mux142(res[13], 1'b0 , W4[13], select[4]);
mux_2_1_helper mux143(res[14], 1'b0 , W4[14], select[4]);
mux_2_1_helper mux144(res[15], 1'b0 , W4[15], select[4]);
mux_2_1_helper mux145(res[16], W4[0] , W4[16], select[4]);
mux_2_1_helper mux146(res[17], W4[1] , W4[17], select[4]);
mux_2_1_helper mux147(res[18], W4[2] , W4[18], select[4]);
mux_2_1_helper mux148(res[19], W4[3] , W4[19], select[4]);
mux_2_1_helper mux149(res[20], W4[4] , W4[20], select[4]);
mux_2_1_helper mux150(res[21], W4[5] , W4[21], select[4]);
mux_2_1_helper mux151(res[22], W4[6] , W4[22], select[4]);
mux_2_1_helper mux152(res[23], W4[7] , W4[23], select[4]);
mux_2_1_helper mux153(res[24], W4[8] , W4[24], select[4]);
mux_2_1_helper mux154(res[25], W4[9] , W4[25], select[4]);
mux_2_1_helper mux155(res[26], W4[10] , W4[26], select[4]);
mux_2_1_helper mux156(res[27], W4[11] , W4[27], select[4]);
mux_2_1_helper mux157(res[28], W4[12] , W4[28], select[4]);
mux_2_1_helper mux158(res[29], W4[13] , W4[29], select[4]);
mux_2_1_helper mux159(res[30], W4[14] , W4[30], select[4]);
mux_2_1_helper mux160(res[31], W4[15] , W4[31], select[4]);

endmodule
 